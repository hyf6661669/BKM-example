library verilog;
use verilog.vl_types.all;
entity barc_tb is
end barc_tb;
